* Active Inverting Gain Subcircuit using LF347 Op-amp

.INC ../components/LF347.cir

* Connections:
*   nIN = Voltage Input
*   nOUT = Voltage Output
*   nPP = Positive Op-amp Power Supply (V+)
*   nNN = Negative Op-amp Power Supply (V-)

* NOTE: The defaults for the params are necessary to prevent LTSpice from
* complaining. It is strongly advised to explicitly declare all parameters.
.SUBCKT Active_Inv_Gain_LF347    nIN nOUT nPP nNN    PARAMS: Ri=1k Rf=1k

R_i nIN nV-	 {Ri}
R_f nV- nOUT {Rf}

X_opamp GND nV- nPP nNN nOUT LF347

.ENDS Active_Inv_Gain_LF347
